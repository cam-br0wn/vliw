module lsu_decode
(

);


endmodule