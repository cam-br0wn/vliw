// Top level of whole design

module vliw ()

endmodule