// execution stage for LSU
// this module is designed to make memory accesses

module lsu_execute
(
    input is_load,
    input zero_ext,
    input rs1,
    input rs2,
    input imm,
    output [31:0] wr_addr,
    output [31:0] rd_addr
);


endmodule