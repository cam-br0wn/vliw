// this module actually performs communication with data mem

module lsu_writeback
(
    
);


endmodule